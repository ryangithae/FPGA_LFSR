`timescale 10ns / 10ps
//////////////////////////////////////////////////////////////////////////////////
// Company: PU
// Engineer: Ryan Githae
// 
// Create Date: 07/08/2025 02:17:45 PM
// Design Name: 
// Module Name: lfsr
// Project Name: Linear Feedback Shift Register
// Target Devices: Basys3 FPGA
// Tool Versions: Vivado 2024.2
// Description: A Pseudorandom Number generator using an LFSR.
// 
// Dependencies: anode.sv
// 
// Revision:5
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lfsr 
   #(
    parameter LFSR_WIDTH = 16,
    parameter CYCLES_PER_SECOND = 100_000_000
    )
    (
    // Create the clock signal and enable for the register
    input clk,
    //input enable,
    
    // Creating customizable parameters for FPGA
    input [4:0] SW, 
        
    // Optional seed value to allow starting from different bits
    //input seed_present,
    //input [LFSR_WIDTH:1] seed,
    
    // Storing the number generated by the LFSR for simulation
    //output [LFSR_WIDTH:1] result,
    
    //Lighting up the seven segments
    output logic [3:0] anode,
    output logic [6:0] cathode,
    output logic dp
    );
    
     localparam int MIN_WIDTH = 3;
     localparam int MAX_WIDTH = 16; 
     localparam int CYCLES = CYCLES_PER_SECOND;
     localparam int COUNTER_WIDTH = $clog2(CYCLES);
    
    // registers to hold the bits(has a default of LFSR_WIDTH'b1) (A non-zero seed is needed to ensure randomness)
    // and the result of the xnor
    reg [LFSR_WIDTH:1] r_LFSR = 16'd5;
    reg xnor_result;
    reg [COUNTER_WIDTH - 1:0] one_second_counter = '0;
    wire enable;
    
    wire [4:0] switch_forced;
    wire [LFSR_WIDTH:1] encoded;
    
    // forcing the LFSR width to be in between 3 and 16 bits for validity
    assign switch_forced = (SW[4:0] < MIN_WIDTH) ? MIN_WIDTH : (SW[4:0] > MAX_WIDTH) ? MAX_WIDTH : SW[4:0];
    
    sevenseg my_display(
        .clk(clk),
        .reset(1'b0),
        .encoded(encoded),
        .decimal_point(dp),
        .anode(anode),
        .cathode(cathode)
        );
     
     // masking logic to handle dynamic sizing of the lenght of the LFSR
     wire [LFSR_WIDTH:1] dynamic_mask;
     genvar i;
     generate
        for (i = 1;i <= LFSR_WIDTH; i = i+1) begin
            assign dynamic_mask[i] = (i <= switch_forced) ? 1'b1 : 1'b0;
        end
     endgenerate
    
    always_ff@(posedge clk) begin
        if(one_second_counter > 99999999) 
            one_second_counter <= '0;
        else
            one_second_counter <= one_second_counter + 1;
     end
     
     assign enable = (one_second_counter == 99999999) ? 1'b1 : 1'b0;
     
    // load the LFSR with the seed value if a pulse is detected
    // otherwise run the LFSR regularly
    always_ff@ (posedge clk) begin    
        //if (enable == 1'b1) begin
           // if (seed_present == 1'b1)
           //     r_LFSR <= seed;
             //else
       if (enable == 1'b1)
            r_LFSR <= ({r_LFSR[LFSR_WIDTH - 1:1], xnor_result} & dynamic_mask);
    end 
    
    
    // combinatinal block of the XNOR assignment of the values
    // Case statements handle where to perform the XNOR "taps" as 
    // recommended by this paper: https://docs.amd.com/v/u/en-US/xapp052
    always_comb begin
     unique case (switch_forced)
        3: begin
            xnor_result = r_LFSR[3] ^~ r_LFSR[2];
        end
        4: begin
            xnor_result = ~(r_LFSR[4] ^ r_LFSR[3]);
        end
        5: begin
             xnor_result = r_LFSR[5] ^~ r_LFSR[3];
        end
        6: begin
            xnor_result = r_LFSR[6] ^~ r_LFSR[5];
        end
        7: begin
            xnor_result = r_LFSR[7] ^~ r_LFSR[6];
        end
        8: begin
            xnor_result = r_LFSR[8] ^~ r_LFSR[6] ^~ r_LFSR[5] ^~ r_LFSR[4];
        end
        9: begin
            xnor_result = r_LFSR[9] ^~ r_LFSR[5];
        end
        10: begin
            xnor_result = r_LFSR[10] ^~ r_LFSR[7];
        end
        11: begin
            xnor_result = r_LFSR[11] ^~ r_LFSR[9];
        end
        12: begin
            xnor_result = r_LFSR[12] ^~ r_LFSR[6] ^~ r_LFSR[4] ^~ r_LFSR[1];
        end
        13: begin
            xnor_result = r_LFSR[13] ^~ r_LFSR[4] ^~ r_LFSR[3] ^~ r_LFSR[1];
        end  
        14: begin
            xnor_result = r_LFSR[14] ^~ r_LFSR[5] ^~ r_LFSR[3] ^~ r_LFSR[1];
        end
        15: begin   
            xnor_result = r_LFSR[15] ^~ r_LFSR[14];
        end
        16: begin
            xnor_result = r_LFSR[16] ^~ r_LFSR[15] ^~ r_LFSR[13] ^~ r_LFSR[4];
        end
        /* 2^16 is the maximum that can be shown on a seven seg display with four segments in hex mode.
        17: begin
            xnor_result = r_LFSR[17] ^~ r_LFSR[14];
        end
        18: begin
            xnor_result = r_LFSR[18] ^~ r_LFSR[11];
        end
        19: begin
            xnor_result = r_LFSR[19] ^~ r_LFSR[6] ^~ r_LFSR[2] ^~ r_LFSR[1];
        end
        20: begin
            xnor_result = r_LFSR[20] ^~ r_LFSR[17];
        end
        21: begin
            xnor_result = r_LFSR[21] ^~ r_LFSR[19];
        end
        22: begin
            xnor_result = r_LFSR[22] ^~ r_LFSR[21];
        end
        23: begin
            xnor_result = r_LFSR[23] ^~ r_LFSR[18];
        end
        24: begin
            xnor_result = r_LFSR[24] ^~ r_LFSR[23] ^~ r_LFSR[22] ^~ r_LFSR[17];
        end
        25: begin
            xnor_result = r_LFSR[25] ^~ r_LFSR[22];
        end
        26: begin
            xnor_result = r_LFSR[26] ^~ r_LFSR[6] ^~ r_LFSR[2] ^~ r_LFSR[1];
        end
        27: begin
             xnor_result = r_LFSR[27] ^~ r_LFSR[5] ^~ r_LFSR[2] ^~ r_LFSR[1];
        end
        28: begin
             xnor_result = r_LFSR[28] ^~ r_LFSR[25];
        end
        29: begin
             xnor_result = r_LFSR[29] ^~ r_LFSR[27];
        end
        30: begin
              xnor_result = r_LFSR[30] ^~ r_LFSR[6] ^~ r_LFSR[4] ^~ r_LFSR[1];
        end
        31: begin
              xnor_result = r_LFSR[31] ^~ r_LFSR[28];
        end
        32: begin
             xnor_result = r_LFSR[32] ^~ r_LFSR[22] ^~ r_LFSR[2] ^~ r_LFSR[1]; 
        end
        */
        default: xnor_result = 1'b0;
    endcase
  end
  
  //assign result = r_LFSR[LFSR_WIDTH:1];
  // assign the LFSR result to the wire that will handle displaying the result
  // on the seven segment display
  assign encoded = r_LFSR;
                
endmodule
